module cacheL2();

endmodule
