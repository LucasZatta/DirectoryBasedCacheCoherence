module processor0();
endmodule
