module processor1();
endmodule
