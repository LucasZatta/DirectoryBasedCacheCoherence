module cacheL1();

endmodule
